// gpio_test_pkg.sv

`include "uvm_macros.svh"

package gpio_test_pkg;

import uvm_pkg::*;

import gpio_env_pkg::*;

`include "gpio_base_test.sv"

endpackage
