// gpio_env_pkg.sv

`include "uvm_macros.svh"

package gpio_env_pkg;

import uvm_pkg::*;

`include "gpio_env_config.sv"
`include "gpio_env.sv"

endpackage
